library verilog;
use verilog.vl_types.all;
entity mux_4to1 is
    port(
        i0              : in     vl_logic_vector(3 downto 0);
        i1              : in     vl_logic_vector(3 downto 0);
        i2              : in     vl_logic_vector(3 downto 0);
        i3              : in     vl_logic_vector(3 downto 0);
        sel             : in     vl_logic_vector(1 downto 0);
        \out\           : out    vl_logic_vector(3 downto 0)
    );
end mux_4to1;
