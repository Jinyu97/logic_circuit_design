library verilog;
use verilog.vl_types.all;
entity or_tb is
end or_tb;
