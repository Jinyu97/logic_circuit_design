library verilog;
use verilog.vl_types.all;
entity cnt_up_down_tb is
end cnt_up_down_tb;
