library verilog;
use verilog.vl_types.all;
entity rcc_tb is
end rcc_tb;
