//??? ??? ?? ???
module SR_latch(Q, Qbar, Sbar, Rbar);

//?? ??
output Q, Qbar;
input Sbar, Rbar;

//Verilog ?????? nand ???? ??
nand n1(Q, Sbar, Qbar);
nand n2(Qbar, Rbar, Q);

endmodule
