module RCC_tb;

reg clk;
reg reset;
wire [3:0] q;

//?? ??? ??
RCC r1(q, clk, reset);

//?? ???? ??? clk ??? ??. ??=10
initial
	clk=1'b0; //clk? 0?? ??
always
	#5 clk = ~clk; //? 5?????? clk ?? ???.
	
//?? ???? ??? reset ??? ??
//reset ??? 0?? 20 ??? 200?? 220?? ???.
initial
begin
	reset = 1'b1;
	#15 reset = 1'b0;
	#180 reset = 1'b1;
	#10 reset = 1'b0;
	#20 $finish; //?????? ??
	end

//??? ??
initial
	$monitor($time, " Output q = %d", q);

endmodule