module OR(Y, A, B);
	input A, B;
	output Y;
	
	or (Y, A, B);
endmodule
