library verilog;
use verilog.vl_types.all;
entity and_tb is
end and_tb;
